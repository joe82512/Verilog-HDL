// ==================== design.sv ====================
// Code your design here

//waveform: Icarus Verilog 0.9.7
//synthesis: Mentor Precision 2021.1+run.do

// 動態(loop次數未知) + 不帶內嵌時序 -> 不可綜合 !!!
module count_ones_c (bit_count, data, clk, reset);
    parameter data_width = 4;
    parameter count_width = 3;
    output [count_width-1: 0] bit_count;
    input  [data_width-1: 0]  data;
    input                     clk, reset;
    reg    [count_width-1: 0] count, bit_count, index;
    reg    [data_width-1: 0]  temp;

    always @ (posedge clk)
        if (reset) begin
            count = 0;
            bit_count = 0;
        end
        else begin
            count = 0;
            temp = data;
            for (index = 0; | temp; index = index + 1) begin //loop次數未知
                if (temp[0] ) count = count + 1;
                temp = temp >> 1;
            end
            bit_count = count;
        end
endmodule

// testcase
module t_count_ones_c ();
    parameter data_width = 4;
    parameter count_width = 3;
    wire [count_width-1:0] bit_count;
    reg  [data_width-1:0]  data;
    reg                    clk, reset;
 
    count_ones_c M0 (bit_count, data, clk, reset);

    //EPWave
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars;
        #500 $finish;
    end

    initial fork
        reset = 1;  // modified 5-17-2002 for longer reset
        #10 reset = 0;
        #200 reset = 1;
        #211 reset = 0;
    join

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    initial begin
        #10 data = 4'hf;
        #40 data = 4'ha;
        #40 data = 4'h5;
        #40 data = 4'hb;
        #40 data = 4'h9;
        #40 data = 4'h0;
        #40 data = 4'hc;
    end
endmodule